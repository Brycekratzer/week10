module top
#(
    parameter DIVIDE_BY = 17 // Use this when passing in to your clock div!
    // The test bench will set it appropriately
)
(
    input [7:0] sw, // A and B
    input clk, // 100 MHz board clock
    input btnC, // Reset
    output [3:0] an, // 7seg anodes
    output [6:0] seg // 7seg segments
);
    wire reset = btnC;
    wire clock = div_clock;

    clock_div #(.DIVIDE_BY(DIVIDE_BY)) clk_div(
        .clock(clk),
        .reset(reset),
        .output(div_clock)
    );

    seven_seg_scanner seven_scnner(
        
    )
    // Instantiate the clock divider...
    // ... wire it up to the scanner
    // ... wire the scanner to the decoder

    // Wire up the math block into the decoder

    // Do not forget to wire up resets!!

endmodule